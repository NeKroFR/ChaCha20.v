`ifndef CHACHA20_DEFS_VH
`define CHACHA20_DEFS_VH

// Constants for ChaCha20
`define CHACHA20_CONST_0 32'h61707865
`define CHACHA20_CONST_1 32'h3320646e
`define CHACHA20_CONST_2 32'h79622d32
`define CHACHA20_CONST_3 32'h6b206574

// Block sizes
`define CHACHA20_BLOCK_SIZE_BITS 512
`define CHACHA20_BLOCK_SIZE_BYTES 64
`define CHACHA20_BLOCK_SIZE_WORDS 16

// Key sizes
`define CHACHA20_KEY_SIZE_BITS 256
`define CHACHA20_KEY_SIZE_BYTES 32
`define CHACHA20_KEY_SIZE_WORDS 8

// Nonce sizes
`define CHACHA20_NONCE_SIZE_BITS 96
`define CHACHA20_NONCE_SIZE_BYTES 12
`define CHACHA20_NONCE_SIZE_WORDS 3

// Counter sizes
`define CHACHA20_COUNTER_SIZE_BITS 32
`define CHACHA20_COUNTER_SIZE_BYTES 4
`define CHACHA20_COUNTER_SIZE_WORDS 1

// Number of rounds
`define CHACHA20_ROUNDS 20

`endif // CHACHA20_DEFS_VH
